module Decoder(a, q);

input [4:0]a;
output reg [31:0]q;

always @ (*)
begin 
	case(a)
	5'b00000: q=32'b0000_0000_0000_0000_0000_0000_0000_0001;
	5'b00001: q=32'b0000_0000_0000_0000_0000_0000_0000_0010;
	5'b00010: q=32'b0000_0000_0000_0000_0000_0000_0000_0100;
	5'b00011: q=32'b0000_0000_0000_0000_0000_0000_0000_1000;
	5'b00100: q=32'b0000_0000_0000_0000_0000_0000_0001_0000;
	5'b00101: q=32'b0000_0000_0000_0000_0000_0000_0010_0000;
	5'b00110: q=32'b0000_0000_0000_0000_0000_0000_0100_0000;
	5'b00111: q=32'b0000_0000_0000_0000_0000_0000_1000_0000;
	5'b01000: q=32'b0000_0000_0000_0000_0000_0001_0000_0000;
	5'b01001: q=32'b0000_0000_0000_0000_0000_0010_0000_0000;
	5'b01010: q=32'b0000_0000_0000_0000_0000_0100_0000_0000;
	5'b01011: q=32'b0000_0000_0000_0000_0000_1000_0000_0000;
	5'b01100: q=32'b0000_0000_0000_0000_0001_0000_0000_0000;
	5'b01101: q=32'b0000_0000_0000_0000_0010_0000_0000_0000;
	5'b01110: q=32'b0000_0000_0000_0000_0100_0000_0000_0000;
	5'b01111: q=32'b0000_0000_0000_0000_1000_0000_0000_0000;
	5'b10000: q=32'b0000_0000_0000_0001_0000_0000_0000_0000;
	5'b10001: q=32'b0000_0000_0000_0010_0000_0000_0000_0000;
	5'b10010: q=32'b0000_0000_0000_0100_0000_0000_0000_0000;
	5'b10011: q=32'b0000_0000_0000_1000_0000_0000_0000_0000;
	5'b10100: q=32'b0000_0000_0001_0000_0000_0000_0000_0000;
	5'b10101: q=32'b0000_0000_0010_0000_0000_0000_0000_0000;
	5'b10110: q=32'b0000_0000_0100_0000_0000_0000_0000_0000;
	5'b10111: q=32'b0000_0000_1000_0000_0000_0000_0000_0000;
	5'b11000: q=32'b0000_0001_0000_0000_0000_0000_0000_0000;
	5'b11001: q=32'b0000_0010_0000_0000_0000_0000_0000_0000;
	5'b11010: q=32'b0000_0100_0000_0000_0000_0000_0000_0000;
	5'b11011: q=32'b0000_1000_0000_0000_0000_0000_0000_0000;
	5'b11100: q=32'b0001_0000_0000_0000_0000_0000_0000_0000;
	5'b11101: q=32'b0010_0000_0000_0000_0000_0000_0000_0000;
	5'b11110: q=32'b0100_0000_0000_0000_0000_0000_0000_0000;
	5'b11111: q=32'b1000_0000_0000_0000_0000_0000_0000_0000;
	endcase
end
endmodule
